//ID/EX�׶εļĴ���
// ʵ��������ִ�н׶�֮��ļĴ�����������׶εĽ������һ��ʱ�����ڴ��ݵ�ִ�н׶�
//////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps
`include "defines.v"

module id_ex(

	input	wire clk,
	input wire rst,

	//���Կ���ģ�����Ϣ
	input wire[5:0]	 stall,
	
	//������׶δ��ݵ���Ϣ
	input wire[`AluOpBus]         id_aluop,//����׶ε�ָ��Ҫ���е����������
	input wire[`AluSelBus]        id_alusel,//����׶ε�ָ��Ҫ���е������������
	input wire[`RegBus]           id_reg1,//����׶ε�ָ��Ҫ���е������Դ������1
	input wire[`RegBus]           id_reg2,//����׶ε�ָ��Ҫ���е������Դ������2?
	input wire[`RegAddrBus]       id_wd,//����׶ε�ָ��Ҫд���Ŀ�ļĴ�����ַ
	input wire                    id_wreg,//����׶ε�ָ���Ƿ���Ҫд���Ŀ�ļĴ���
	input wire[`RegBus]           id_link_address,//��ǰ��������׶ε�ָ���Ƿ�λ���ӳٲ�
	input wire                    id_is_in_delayslot,//��������׶ε�ת��ָ��Ҫ����ķ��ص�ַ
	input wire                    next_inst_in_delayslot_i,	//��һ����������׶ε�ָ���Ƿ�λ���ӳٲ�	
	
	//���ݵ�ִ�н׶ε���Ϣ
	output reg[`AluOpBus]         ex_aluop,//ִ�н׶ε�ָ��Ҫ���е����������
	output reg[`AluSelBus]        ex_alusel,//ִ�н׶ε�ָ��Ҫ���е������������
	output reg[`RegBus]           ex_reg1,//ִ�н׶ε�ָ��Ҫ���е������Դ������1
	output reg[`RegBus]           ex_reg2,//ִ�н׶ε�ָ��Ҫ���е������Դ������2
	output reg[`RegAddrBus]       ex_wd,//ִ�н׶ε�ָ��Ҫд���Ŀ�ļĴ�����ַ
	output reg                    ex_wreg,//ִ�н׶ε�ָ���Ƿ���Ҫд���Ŀ�ļĴ���
	output reg[`RegBus]           ex_link_address,//����ִ�н׶ε�ת��ָ��Ҫ����ķ��ص�ַ
  output reg                    ex_is_in_delayslot,//��ǰ����ִ�н׶ε�ָ���Ƿ�λ���ӳٲ�
	output reg                    is_in_delayslot_o	//��ǰ��������׶ε�ָ���Ƿ�λ���ӳٲ�
	
);

	always @ (posedge clk) begin
		if (rst == `RstEnable) begin
			ex_aluop <= `EXE_NOP_OP;
			ex_alusel <= `EXE_RES_NOP;
			ex_reg1 <= `ZeroWord;
			ex_reg2 <= `ZeroWord;
			ex_wd <= `NOPRegAddr;
			ex_wreg <= `WriteDisable;
			ex_link_address <= `ZeroWord;
			ex_is_in_delayslot <= `NotInDelaySlot;
	    is_in_delayslot_o <= `NotInDelaySlot;			
	    
	    //1���� stall��2��Ϊ Stop��stall��3��ΪNoStopʱ����ʾ����׶���ͣ��
	    //��ִ�н׶μ���������ʹ�ÿ�ָ����Ϊ��һ�����ڽ���ִ�н׶ε�ָ��
	    //2����stall��2��ΪNoStop ʱ������׶μ�����������ָ�����ִ�н׶�
	    //3����������£�����ִ�н׶εļĴ���ex aluop��
	    //ex_alusel��ex_reg1��?ex_reg2��ex _wd��ex_wreg ���䡤
	  
		end else if(stall[2] == `Stop && stall[3] == `NoStop) begin
			ex_aluop <= `EXE_NOP_OP;
			ex_alusel <= `EXE_RES_NOP;
			ex_reg1 <= `ZeroWord;
			ex_reg2 <= `ZeroWord;
			ex_wd <= `NOPRegAddr;
			ex_wreg <= `WriteDisable;	
			ex_link_address <= `ZeroWord;
	    ex_is_in_delayslot <= `NotInDelaySlot;			
	    
	//����ˮ������׶�û�б���ͣʱ��ID/EXģ����ʱ�������ؽ������ӵ����봫�ݵ���Ӧ�����    
		end else if(stall[2] == `NoStop) begin		
			ex_aluop <= id_aluop;
			ex_alusel <= id_alusel;
			ex_reg1 <= id_reg1;
			ex_reg2 <= id_reg2;
			ex_wd <= id_wd;
			ex_wreg <= id_wreg;		
			
			
			ex_link_address <= id_link_address;
			ex_is_in_delayslot <= id_is_in_delayslot;
	    is_in_delayslot_o <= next_inst_in_delayslot_i;				
		end
	end
	
endmodule